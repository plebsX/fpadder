module fpadder
(
	output	logic [31:0] sum,
	output	logic ready,
	input	logic [31:0] a,
	input	logic clock,
	input	logic nreset
);
//enum {start,loada, loadb,sign,exp_equal,add_m,normalise} present_state, next_state;
enum {start,loada,loadb,zerock,exp_equal,add_m,normalise} present_state, next_state;
logic	[25:0]	mx;
logic	[25:0]	my;
logic 	[25:0]	m_result;

logic	[7:0]	ex;
logic	[7:0]	ey;
logic 	[7:0]	e_result;

logic 	[31:0]	ix;
logic	[31:0]	iy;
logic	[31:0]  result;

//assign result=(present_state==start)?{m_result[25],e_result[7:0],m_result[22:0]}:'b0;
assign sum = (present_state==start)?{m_result[25],e_result[7:0],m_result[22:0]}:'bX;
assign ready = (present_state==start)? 1:0;
//always_ff @(posedge clock or negedge nreset) begin
//	if(nreset == 1'b0)begin
//		sum <= 'b0;
//	end
//	else begin
//		if(present_state == start)
//		begin
//			sum <= {m_result[25],e_result[7:0],m_result[22:0]};
//		end
//		else
//			sum <= sum;
//	end
//end

//always_ff @(posedge clock or negedge nreset) begin
//	if(nreset == 1'b0)begin
//		ready <= 'b0;
//	end
//	else begin
//		if(present_state == start)
//		begin
//			ready <= 1'b1;
//		end
//		else
//			ready <= 1'b0;
//	end
//end

always_ff  @(posedge clock or negedge nreset)begin
    if(nreset==1'b0)begin
		present_state <= start;
    end
    else begin
		present_state <= next_state;
    end
end

always_comb
begin
	unique case(present_state)
		start:begin
			next_state = loada;
		end
		loada:begin
			ix = a;
			ex = a[30:23];
			mx = {a[31],1'b0,1'b1,a[22:0]};
			next_state = loadb;
		end
		loadb:begin
			iy = a;
			ey = a[30:23];
			my = {a[31],1'b0,1'b1,a[22:0]};
			next_state = zerock;
		end
		zerock:begin
			if(ix == 0)
			begin
				{e_result, m_result} = {ey,my};
				next_state = start;
			end	
			else if(iy==0)
			begin
				{e_result, m_result} = {ex,mx};
				next_state = start;

			end
			else
				next_state = exp_equal;
		end
		exp_equal:begin
			if(ex == ey)
			begin
				e_result = ex;
				next_state = add_m;
			end
			else if(ex > ey)
			begin
				ey = ey + 1;
				my[24:0] = {1'b0,my[24:1]};
				if(my == 0)
				begin
					m_result = mx;
					e_result = ex;
					next_state = start;
				end
				else
					next_state = exp_equal;	
			end
			else if(ex < ey)
			begin
				ex = ex + 1;
				mx[24:0] <= {1'b0,mx[24:1]};
				if(mx == 0)
				begin
					m_result = my;
					e_result = ey;
					next_state = start;
				end
				else
					next_state = exp_equal;
			end
		end
		add_m : begin
			if((mx[25] == my[25]))
			begin
				m_result[25] = mx[25];
				m_result[24:0] = mx[24:0]+my[24:0];
			end
			else
			begin
				if(mx[24:0]>my[24:0])//mx > my
				begin
					m_result[25] = mx[25];
					m_result[24:0] = mx[24:0] - my[24:0];
				end
				else
				begin
					m_result[25] = my[25];
					m_result[24:0] = my[24:0] - mx[24:0];
				end
			end
			next_state = normalise;	
		
		end
		normalise:begin
			if(m_result[24]==1)
			begin
				m_result[24:0] = {1'b0,m_result[24:1]};
				e_result = e_result +1;
				next_state = start;
			end
			else if(m_result[23]==0)
			begin
				m_result = {m_result[23:0],1'b0};
				e_result = e_result -1;
				next_state = normalise;
			end
			else
				next_state = start;
		end
	endcase
end


endmodule





















